`ifndef __AXI_ADDRESSES__
`define __AXI_ADDRESSES__

`define KEY_ADDR  32'h00000100
`define DATA_ADDR 32'h00000200
`define ADDR_MASK 32'hFFFFF000

`endif
